module req_gen (clk, rst, out_ptr, out_ptr_vld);

input clk;
input rst;
output out_ptr_vld;
output [7:0] out_ptr;

wire vdd = 1'b1;
wire gnd = 1'b0;

INVX4 INVX4_1 ( .A(_14_), .Y(_15_) );
NOR2X1 NOR2X1_1 ( .A(_0__5_), .B(_0__4_), .Y(_16_) );
NOR2X1 NOR2X1_2 ( .A(_0__7_), .B(_0__6_), .Y(_17_) );
AND2X2 AND2X2_1 ( .A(_16_), .B(_17_), .Y(_18_) );
INVX1 INVX1_1 ( .A(_0__3_), .Y(_19_) );
NOR2X1 NOR2X1_3 ( .A(_0__2_), .B(_19_), .Y(_20_) );
NAND3X1 NAND3X1_1 ( .A(_0__0_), .B(_20_), .C(_18_), .Y(_21_) );
NAND3X1 NAND3X1_2 ( .A(_0__1_), .B(_0__3_), .C(_0__2_), .Y(_22_) );
INVX1 INVX1_2 ( .A(_22_), .Y(_23_) );
NAND2X1 NAND2X1_1 ( .A(_23_), .B(_18_), .Y(_24_) );
AND2X2 AND2X2_2 ( .A(_0__3_), .B(_0__2_), .Y(_25_) );
INVX1 INVX1_3 ( .A(_0__0_), .Y(_26_) );
NOR2X1 NOR2X1_4 ( .A(_0__1_), .B(_26_), .Y(_27_) );
NAND3X1 NAND3X1_3 ( .A(_25_), .B(_27_), .C(_18_), .Y(_28_) );
NAND3X1 NAND3X1_4 ( .A(_24_), .B(_21_), .C(_28_), .Y(_29_) );
NOR2X1 NOR2X1_5 ( .A(_0__3_), .B(_0__2_), .Y(_30_) );
NOR2X1 NOR2X1_6 ( .A(_0__0_), .B(_30_), .Y(_31_) );
NAND3X1 NAND3X1_5 ( .A(_22_), .B(_31_), .C(_18_), .Y(_32_) );
INVX1 INVX1_4 ( .A(_0__1_), .Y(_33_) );
NOR2X1 NOR2X1_7 ( .A(_0__0_), .B(_33_), .Y(_34_) );
NAND3X1 NAND3X1_6 ( .A(_34_), .B(_30_), .C(_18_), .Y(_35_) );
NAND2X1 NAND2X1_2 ( .A(_0__0_), .B(_0__1_), .Y(_36_) );
NOR3X1 NOR3X1_1 ( .A(_0__3_), .B(_0__2_), .C(_36_), .Y(_37_) );
INVX1 INVX1_5 ( .A(_0__2_), .Y(_38_) );
NOR3X1 NOR3X1_2 ( .A(_0__3_), .B(_26_), .C(_38_), .Y(_39_) );
OAI21X1 OAI21X1_1 ( .A(_37_), .B(_39_), .C(_18_), .Y(_40_) );
NAND3X1 NAND3X1_7 ( .A(_32_), .B(_35_), .C(_40_), .Y(_41_) );
AND2X2 AND2X2_3 ( .A(_18_), .B(_20_), .Y(_42_) );
INVX1 INVX1_6 ( .A(_36_), .Y(_43_) );
NAND2X1 NAND2X1_3 ( .A(_16_), .B(_17_), .Y(_44_) );
NAND3X1 NAND3X1_8 ( .A(_26_), .B(_0__1_), .C(_25_), .Y(_45_) );
NAND3X1 NAND3X1_9 ( .A(_0__0_), .B(_0__2_), .C(_19_), .Y(_46_) );
AOI21X1 AOI21X1_1 ( .A(_45_), .B(_46_), .C(_44_), .Y(_47_) );
AOI21X1 AOI21X1_2 ( .A(_42_), .B(_43_), .C(_47_), .Y(_48_) );
OAI21X1 OAI21X1_2 ( .A(_29_), .B(_41_), .C(_48_), .Y(_49_) );
AOI22X1 AOI22X1_1 ( .A(i_ptr_seq_gen_start_0_), .B(_15_), .C(_1_), .D(_49_), .Y(_50_) );
INVX1 INVX1_7 ( .A(_50_), .Y(i_ptr_seq_gen_cur_0_) );
NAND2X1 NAND2X1_4 ( .A(_0__3_), .B(_0__2_), .Y(_51_) );
NOR3X1 NOR3X1_3 ( .A(_0__0_), .B(_33_), .C(_51_), .Y(_52_) );
NAND2X1 NAND2X1_5 ( .A(_52_), .B(_18_), .Y(_53_) );
NAND3X1 NAND3X1_10 ( .A(_20_), .B(_27_), .C(_18_), .Y(_54_) );
NAND3X1 NAND3X1_11 ( .A(_53_), .B(_54_), .C(_40_), .Y(_55_) );
AOI22X1 AOI22X1_2 ( .A(i_ptr_seq_gen_start_1_), .B(_15_), .C(_1_), .D(_55_), .Y(_56_) );
INVX1 INVX1_8 ( .A(_56_), .Y(i_ptr_seq_gen_cur_1_) );
INVX1 INVX1_9 ( .A(i_ptr_seq_gen_start_2_), .Y(_57_) );
NOR2X1 NOR2X1_8 ( .A(_29_), .B(_41_), .Y(_58_) );
NAND3X1 NAND3X1_12 ( .A(_0__1_), .B(_39_), .C(_18_), .Y(_59_) );
AND2X2 AND2X2_4 ( .A(_59_), .B(_21_), .Y(_60_) );
NAND3X1 NAND3X1_13 ( .A(_28_), .B(_35_), .C(_60_), .Y(_61_) );
OAI21X1 OAI21X1_3 ( .A(_61_), .B(_58_), .C(_1_), .Y(_62_) );
OAI21X1 OAI21X1_4 ( .A(_57_), .B(_14_), .C(_62_), .Y(i_ptr_seq_gen_cur_2_) );
INVX1 INVX1_10 ( .A(i_ptr_seq_gen_start_3_), .Y(_63_) );
INVX1 INVX1_11 ( .A(_37_), .Y(_64_) );
OAI21X1 OAI21X1_5 ( .A(_44_), .B(_64_), .C(_59_), .Y(_65_) );
OAI21X1 OAI21X1_6 ( .A(_65_), .B(_29_), .C(_1_), .Y(_66_) );
OAI21X1 OAI21X1_7 ( .A(_63_), .B(_14_), .C(_66_), .Y(i_ptr_seq_gen_cur_3_) );
AND2X2 AND2X2_5 ( .A(_15_), .B(gnd), .Y(i_ptr_seq_gen_cur_4_) );
AND2X2 AND2X2_6 ( .A(_15_), .B(gnd), .Y(i_ptr_seq_gen_cur_5_) );
AND2X2 AND2X2_7 ( .A(_15_), .B(gnd), .Y(i_ptr_seq_gen_cur_6_) );
AND2X2 AND2X2_8 ( .A(_15_), .B(gnd), .Y(i_ptr_seq_gen_cur_7_) );
NOR2X1 NOR2X1_9 ( .A(_46_), .B(_44_), .Y(_67_) );
NAND3X1 NAND3X1_14 ( .A(_21_), .B(_28_), .C(_35_), .Y(_68_) );
AOI21X1 AOI21X1_3 ( .A(_0__1_), .B(_67_), .C(_68_), .Y(_69_) );
OAI21X1 OAI21X1_8 ( .A(_29_), .B(_41_), .C(_69_), .Y(_70_) );
AOI22X1 AOI22X1_3 ( .A(i_ptr_seq_gen_start_2_), .B(_15_), .C(_1_), .D(_70_), .Y(_71_) );
OAI21X1 OAI21X1_9 ( .A(gnd), .B(gnd), .C(_15_), .Y(_72_) );
OAI21X1 OAI21X1_10 ( .A(gnd), .B(gnd), .C(_15_), .Y(_73_) );
AND2X2 AND2X2_9 ( .A(_72_), .B(_73_), .Y(_2_) );
NAND2X1 NAND2X1_6 ( .A(_2_), .B(_56_), .Y(_3_) );
NOR2X1 NOR2X1_10 ( .A(_3_), .B(i_ptr_seq_gen_cur_3_), .Y(_4_) );
NAND3X1 NAND3X1_15 ( .A(_50_), .B(_4_), .C(_71_), .Y(i_ptr_seq_gen_cur_vld) );
AND2X2 AND2X2_10 ( .A(_27_), .B(_25_), .Y(_5_) );
OAI21X1 OAI21X1_11 ( .A(_23_), .B(_5_), .C(_18_), .Y(_7_) );
AOI22X1 AOI22X1_4 ( .A(_18_), .B(_37_), .C(_0__1_), .D(_67_), .Y(_8_) );
NAND3X1 NAND3X1_16 ( .A(_21_), .B(_7_), .C(_8_), .Y(_9_) );
AOI22X1 AOI22X1_5 ( .A(i_ptr_seq_gen_start_3_), .B(_15_), .C(_1_), .D(_9_), .Y(_10_) );
AND2X2 AND2X2_11 ( .A(_56_), .B(_2_), .Y(_11_) );
NAND3X1 NAND3X1_17 ( .A(_10_), .B(_11_), .C(_50_), .Y(_12_) );
NOR2X1 NOR2X1_11 ( .A(i_ptr_seq_gen_cur_2_), .B(_12_), .Y(i_ptr_seq_gen_start_rdy) );
INVX1 INVX1_12 ( .A(rst), .Y(_6_) );
DFFPOSX1 DFFPOSX1_1 ( .CLK(clk), .D(i_ptr_seq_gen_cur_0_), .Q(_0__0_) );
DFFPOSX1 DFFPOSX1_2 ( .CLK(clk), .D(i_ptr_seq_gen_cur_1_), .Q(_0__1_) );
DFFPOSX1 DFFPOSX1_3 ( .CLK(clk), .D(i_ptr_seq_gen_cur_2_), .Q(_0__2_) );
DFFPOSX1 DFFPOSX1_4 ( .CLK(clk), .D(i_ptr_seq_gen_cur_3_), .Q(_0__3_) );
DFFPOSX1 DFFPOSX1_5 ( .CLK(clk), .D(i_ptr_seq_gen_cur_4_), .Q(_0__4_) );
DFFPOSX1 DFFPOSX1_6 ( .CLK(clk), .D(i_ptr_seq_gen_cur_5_), .Q(_0__5_) );
DFFPOSX1 DFFPOSX1_7 ( .CLK(clk), .D(i_ptr_seq_gen_cur_6_), .Q(_0__6_) );
DFFPOSX1 DFFPOSX1_8 ( .CLK(clk), .D(i_ptr_seq_gen_cur_7_), .Q(_0__7_) );
DFFSR DFFSR_1 ( .CLK(clk), .D(i_ptr_seq_gen_cur_vld), .Q(_1_), .R(_6_), .S(vdd) );
INVX2 INVX2_1 ( .A(i_start_req_gen_n_req_2_), .Y(_75_) );
NOR2X1 NOR2X1_12 ( .A(i_start_req_gen_n_req_1_), .B(i_start_req_gen_n_req_0_), .Y(_76_) );
NAND3X1 NAND3X1_18 ( .A(_75_), .B(i_start_req_gen_n_req_3_), .C(_76_), .Y(i_ptr_seq_gen_start_vld) );
XOR2X1 XOR2X1_1 ( .A(i_start_req_gen_n_req_0_), .B(i_ptr_seq_gen_start_rdy), .Y(_74__0_) );
OR2X2 OR2X2_1 ( .A(i_start_req_gen_n_req_1_), .B(i_ptr_seq_gen_start_rdy), .Y(_77_) );
AND2X2 AND2X2_12 ( .A(i_start_req_gen_n_req_1_), .B(i_start_req_gen_n_req_0_), .Y(_78_) );
OAI21X1 OAI21X1_12 ( .A(_76_), .B(_78_), .C(i_ptr_seq_gen_start_rdy), .Y(_79_) );
AND2X2 AND2X2_13 ( .A(_79_), .B(_77_), .Y(_74__1_) );
NAND3X1 NAND3X1_19 ( .A(i_start_req_gen_n_req_1_), .B(i_start_req_gen_n_req_0_), .C(i_ptr_seq_gen_start_rdy), .Y(_80_) );
XNOR2X1 XNOR2X1_1 ( .A(_80_), .B(i_start_req_gen_n_req_2_), .Y(_74__2_) );
OAI21X1 OAI21X1_13 ( .A(_75_), .B(_80_), .C(i_start_req_gen_n_req_3_), .Y(_81_) );
INVX1 INVX1_13 ( .A(i_start_req_gen_n_req_3_), .Y(_82_) );
INVX1 INVX1_14 ( .A(_80_), .Y(_83_) );
NAND3X1 NAND3X1_20 ( .A(i_start_req_gen_n_req_2_), .B(_82_), .C(_83_), .Y(_84_) );
NAND2X1 NAND2X1_7 ( .A(_81_), .B(_84_), .Y(_74__3_) );
OAI21X1 OAI21X1_14 ( .A(i_start_req_gen_n_req_1_), .B(i_start_req_gen_n_req_0_), .C(i_start_req_gen_n_req_2_), .Y(_85_) );
OAI21X1 OAI21X1_15 ( .A(_76_), .B(_78_), .C(_75_), .Y(_87_) );
NAND3X1 NAND3X1_21 ( .A(_82_), .B(_85_), .C(_87_), .Y(i_ptr_seq_gen_start_0_) );
NAND2X1 NAND2X1_8 ( .A(_75_), .B(_82_), .Y(_88_) );
NOR2X1 NOR2X1_13 ( .A(_78_), .B(_88_), .Y(i_ptr_seq_gen_start_1_) );
NOR2X1 NOR2X1_14 ( .A(i_start_req_gen_n_req_1_), .B(_88_), .Y(i_ptr_seq_gen_start_2_) );
OAI21X1 OAI21X1_16 ( .A(_75_), .B(_76_), .C(_82_), .Y(i_ptr_seq_gen_start_3_) );
INVX2 INVX2_2 ( .A(rst), .Y(_86_) );
DFFSR DFFSR_2 ( .CLK(clk), .D(_74__0_), .Q(i_start_req_gen_n_req_0_), .R(_86_), .S(vdd) );
DFFSR DFFSR_3 ( .CLK(clk), .D(_74__1_), .Q(i_start_req_gen_n_req_1_), .R(_86_), .S(vdd) );
DFFSR DFFSR_4 ( .CLK(clk), .D(_74__2_), .Q(i_start_req_gen_n_req_2_), .R(_86_), .S(vdd) );
DFFSR DFFSR_5 ( .CLK(clk), .D(_74__3_), .Q(i_start_req_gen_n_req_3_), .R(_86_), .S(vdd) );
BUFX2 BUFX2_1 ( .A(_0__0_), .Y(out_ptr[0]) );
BUFX2 BUFX2_2 ( .A(_0__1_), .Y(out_ptr[1]) );
BUFX2 BUFX2_3 ( .A(_0__2_), .Y(out_ptr[2]) );
BUFX2 BUFX2_4 ( .A(_0__3_), .Y(out_ptr[3]) );
BUFX2 BUFX2_5 ( .A(_0__4_), .Y(out_ptr[4]) );
BUFX2 BUFX2_6 ( .A(_0__5_), .Y(out_ptr[5]) );
BUFX2 BUFX2_7 ( .A(_0__6_), .Y(out_ptr[6]) );
BUFX2 BUFX2_8 ( .A(_0__7_), .Y(out_ptr[7]) );
BUFX2 BUFX2_9 ( .A(_1_), .Y(out_ptr_vld) );
INVX1 INVX1_15 ( .A(_1_), .Y(_13_) );
NAND2X1 NAND2X1_9 ( .A(i_ptr_seq_gen_start_vld), .B(_13_), .Y(_14_) );
endmodule
